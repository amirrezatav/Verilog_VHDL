module (o);

endmodule