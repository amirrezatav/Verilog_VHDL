library verilog;
use verilog.vl_types.all;
entity SubtractorTest is
end SubtractorTest;
