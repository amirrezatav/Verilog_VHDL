library verilog;
use verilog.vl_types.all;
entity TOP is
    generic(
        Delay           : integer := 10
    );
end TOP;
