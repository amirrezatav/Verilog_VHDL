module ALU(
    input wire[1:2] sel,
    
);
    
endmodule